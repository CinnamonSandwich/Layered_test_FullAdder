`timescale 1ns / 1ps

interface intf();
  
  logic a;
  logic b;
  logic cin;
  logic sum;
  logic cout;
  
endinterface
